`include "rtl/CPU.v"
`include "rtl/Memory.v"

module Top (
    output something
);
  
endmodule