`include "rtl/Defines.v"

module ALUCtrl (
    input [2:0]  funct3,
    input [6:0]  funct7,
    input [1:0]  aluCtrlOp,
    output reg [3:0] aluOp
);
    always @(*) begin
      case(aluCtrlOp)
        2'b00:  aluOp <= `ALU_OP_ADD;           // Load/Store
        2'b10:  aluOp <= {funct7[5], funct3};   // normal ALUI/ALUR
        2'b01:  case(funct3)                    // bxx
          `BEQ_FUNCT3:  aluOp <= `ALU_OP_EQ;
          `BNE_FUNCT3:  aluOp <= `ALU_OP_NEQ;
          `BLT_FUNCT3:  aluOp <= `ALU_OP_SLT;
          `BGE_FUNCT3:  aluOp <= `ALU_OP_GE;
          `BLTU_FUNCT3: aluOp <= `ALU_OP_SLTU;
          `BGEU_FUNCT3: aluOp <= `ALU_OP_GEU;
          default:      aluOp <= `ALU_OP_XXX;
        endcase
        default: aluOp <= `ALU_OP_XXX;
      endcase
    end
endmodule